module AHBlite_Decoder
#(
    /*RAMCODE enable parameter*/
    parameter Port0_en = 1,
    /************************/

    /*RAMDATA enable parameter*/
    parameter Port1_en = 1,
    /************************/

    /*WaterLight enable parameter*/
    parameter Port2_en = 0,
    /************************/

    /*UART enable parameter*/
    parameter Port3_en=0,
    /************************/

    /*GPIO enable parameter*/
    parameter Port4_en=0,
    /************************/

    /*MicroCode_controller enable parameter*/
    parameter Port5_en = 1,
    /************************/

    /*MicroCode_RAM enable parameter*/
    parameter Port6_en = 1
    /************************/
)(
    input [31:0] HADDR,

    /*RAMCODE OUTPUT SELECTION SIGNAL*/
    output wire P0_HSEL,

    /*WaterLight OUTPUT SELECTION SIGNAL*/
    output wire P1_HSEL,

    /*RAMDATA OUTPUT SELECTION SIGNAL*/
    output wire P2_HSEL,

    /*UART OUTPUT SELECTION SIGNAL*/
    output wire P3_HSEL,       

    /*GPIO OUTPUT SELECTION SIGNAL*/
    output wire P4_HSEL,

    /*MicroCode_controller OUTPUT SELECTION SIGNAL*/
    output wire P5_HSEL,

    /*MicroCode_RAM OUTPUT SELECTION SIGNAL*/
    output wire P6_HSEL      
);

//RAMCODE-----------------------------------

//0x00000000-0x0000ffff
/*Insert RAMCODE decoder code there*/
assign P0_HSEL = (HADDR[31:16] == 16'h0000) ? Port0_en : 1'd0;
/***********************************/



//PERIPHRAL-----------------------------

//0X40000000 WaterLight MODE
//0x40000004 WaterLight SPEED
/*Insert WaterLight decoder code there*/
assign P2_HSEL = 1'd0;
/***********************************/

//0X40000010 UART RX DATA
//0X40000014 UART TX STATE
//0X40000018 UART TX DATA
/*Insert UART decoder code there*/
assign P3_HSEL = 1'b0;
/***********************************/

//0x40000028 OUT  ENABLE
//0X40000024 IN DATA
//0X40000020 OUT DATA
/*Insert GPIO decoder code there*/
assign P4_HSEL = 1'd0;
/***********************************/

//0x40000030 START ADDR
//0X40000034 END ADDR
//0X40000038 ENABLE
//0X4000003c GPIO INPUT (read only)
/*Insert MicroCode_controller decoder code there*/
assign P5_HSEL = (HADDR[31:4] == 28'h4000003) ? Port5_en : 1'd0;
/***********************************/

//0x40001000-0x400013ff
/*Insert MicroCode_controller decoder code there*/
assign P6_HSEL = (HADDR[31:12] == 20'h40001) ? Port6_en : 1'd0;
/***********************************/


//RAMDATA-----------------------------
//0X20000000-0X2000FFFF
/*Insert RAMDATA decoder code there*/
assign P1_HSEL = (HADDR[31:16] == 16'h2000) ? Port1_en : 1'b0;
/***********************************/

endmodule